----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 04/22/2022 10:16:58 PM
-- Design Name: 
-- Module Name: ROM - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.numeric_std.ALL;
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity ROM is
    Port ( addr : in STD_LOGIC_VECTOR (39 downto 0);
           Cout : out STD_LOGIC_VECTOR (19 downto 0));
end ROM;

architecture Behavioral of ROM is
type vector is Array(0 to 1400) of Std_logic_vector(19 downto 0);
Constant memory: vector:=
(0=>x"00000",
1=>x"00000",
2=>x"00000",
3=>x"00000",
4=>x"00000",
5=>x"00000",
6=>x"00000",
7=>x"00000",
8=>x"00000",
9=>x"00000",
10=>x"00000",
11=>x"00000",
12=>x"00000",
13=>x"00000",
14=>x"00001",
15=>x"00001",
16=>x"00001",
17=>x"00001",
18=>x"00001",
19=>x"00001",
20=>x"00001",
21=>x"00001",
22=>x"00001",
23=>x"00001",
24=>x"00001",
25=>x"00001",
26=>x"00001",
27=>x"00001",
28=>x"00002",
29=>x"00002",
30=>x"00002",
31=>x"00002",
32=>x"00002",
33=>x"00002",
34=>x"00002",
35=>x"00002",
36=>x"00002",
37=>x"00002",
38=>x"00002",
39=>x"00002",
40=>x"00002",
41=>x"00002",
42=>x"00003",
43=>x"00003",
44=>x"00003",
45=>x"00003",
46=>x"00003",
47=>x"00003",
48=>x"00003",
49=>x"00003",
50=>x"00003",
51=>x"00003",
52=>x"00003",
53=>x"00003",
54=>x"00003",
55=>x"00003",
56=>x"00004",
57=>x"00004",
58=>x"00004",
59=>x"00004",
60=>x"00004",
61=>x"00004",
62=>x"00004",
63=>x"00004",
64=>x"00004",
65=>x"00004",
66=>x"00004",
67=>x"00004",
68=>x"00004",
69=>x"00004",
70=>x"00005",
71=>x"00005",
72=>x"00005",
73=>x"00005",
74=>x"00005",
75=>x"00005",
76=>x"00005",
77=>x"00005",
78=>x"00005",
79=>x"00005",
80=>x"00005",
81=>x"00005",
82=>x"00005",
83=>x"00005",
84=>x"00006",
85=>x"00006",
86=>x"00006",
87=>x"00006",
88=>x"00006",
89=>x"00006",
90=>x"00006",
91=>x"00006",
92=>x"00006",
93=>x"00006",
94=>x"00006",
95=>x"00006",
96=>x"00006",
97=>x"00006",
98=>x"00007",
99=>x"00007",
100=>x"00007",
101=>x"00007",
102=>x"00007",
103=>x"00007",
104=>x"00007",
105=>x"00007",
106=>x"00007",
107=>x"00007",
108=>x"00007",
109=>x"00007",
110=>x"00007",
111=>x"00007",
112=>x"00008",
113=>x"00008",
114=>x"00008",
115=>x"00008",
116=>x"00008",
117=>x"00008",
118=>x"00008",
119=>x"00008",
120=>x"00008",
121=>x"00008",
122=>x"00008",
123=>x"00008",
124=>x"00008",
125=>x"00008",
126=>x"00009",
127=>x"00009",
128=>x"00009",
129=>x"00009",
130=>x"00009",
131=>x"00009",
132=>x"00009",
133=>x"00009",
134=>x"00009",
135=>x"00009",
136=>x"00009",
137=>x"00009",
138=>x"00009",
139=>x"00009",
140=>x"0000a",
141=>x"0000a",
142=>x"0000a",
143=>x"0000a",
144=>x"0000a",
145=>x"0000a",
146=>x"0000a",
147=>x"0000a",
148=>x"0000a",
149=>x"0000a",
150=>x"0000a",
151=>x"0000a",
152=>x"0000a",
153=>x"0000a",
154=>x"0000b",
155=>x"0000b",
156=>x"0000b",
157=>x"0000b",
158=>x"0000b",
159=>x"0000b",
160=>x"0000b",
161=>x"0000b",
162=>x"0000b",
163=>x"0000b",
164=>x"0000b",
165=>x"0000b",
166=>x"0000b",
167=>x"0000b",
168=>x"0000c",
169=>x"0000c",
170=>x"0000c",
171=>x"0000c",
172=>x"0000c",
173=>x"0000c",
174=>x"0000c",
175=>x"0000c",
176=>x"0000c",
177=>x"0000c",
178=>x"0000c",
179=>x"0000c",
180=>x"0000c",
181=>x"0000c",
182=>x"0000d",
183=>x"0000d",
184=>x"0000d",
185=>x"0000d",
186=>x"0000d",
187=>x"0000d",
188=>x"0000d",
189=>x"0000d",
190=>x"0000d",
191=>x"0000d",
192=>x"0000d",
193=>x"0000d",
194=>x"0000d",
195=>x"0000d",
196=>x"0000e",
197=>x"0000e",
198=>x"0000e",
199=>x"0000e",
200=>x"0000e",
201=>x"0000e",
202=>x"0000e",
203=>x"0000e",
204=>x"0000e",
205=>x"0000e",
206=>x"0000e",
207=>x"0000e",
208=>x"0000e",
209=>x"0000e",
210=>x"0000f",
211=>x"0000f",
212=>x"0000f",
213=>x"0000f",
214=>x"0000f",
215=>x"0000f",
216=>x"0000f",
217=>x"0000f",
218=>x"0000f",
219=>x"0000f",
220=>x"0000f",
221=>x"0000f",
222=>x"0000f",
223=>x"0000f",
224=>x"00010",
225=>x"00010",
226=>x"00010",
227=>x"00010",
228=>x"00010",
229=>x"00010",
230=>x"00010",
231=>x"00010",
232=>x"00010",
233=>x"00010",
234=>x"00010",
235=>x"00010",
236=>x"00010",
237=>x"00010",
238=>x"00011",
239=>x"00011",
240=>x"00011",
241=>x"00011",
242=>x"00011",
243=>x"00011",
244=>x"00011",
245=>x"00011",
246=>x"00011",
247=>x"00011",
248=>x"00011",
249=>x"00011",
250=>x"00011",
251=>x"00011",
252=>x"00012",
253=>x"00012",
254=>x"00012",
255=>x"00012",
256=>x"00012",
257=>x"00012",
258=>x"00012",
259=>x"00012",
260=>x"00012",
261=>x"00012",
262=>x"00012",
263=>x"00012",
264=>x"00012",
265=>x"00012",
266=>x"00013",
267=>x"00013",
268=>x"00013",
269=>x"00013",
270=>x"00013",
271=>x"00013",
272=>x"00013",
273=>x"00013",
274=>x"00013",
275=>x"00013",
276=>x"00013",
277=>x"00013",
278=>x"00013",
279=>x"00013",
280=>x"00014",
281=>x"00014",
282=>x"00014",
283=>x"00014",
284=>x"00014",
285=>x"00014",
286=>x"00014",
287=>x"00014",
288=>x"00014",
289=>x"00014",
290=>x"00014",
291=>x"00014",
292=>x"00014",
293=>x"00014",
294=>x"00015",
295=>x"00015",
296=>x"00015",
297=>x"00015",
298=>x"00015",
299=>x"00015",
300=>x"00015",
301=>x"00015",
302=>x"00015",
303=>x"00015",
304=>x"00015",
305=>x"00015",
306=>x"00015",
307=>x"00015",
308=>x"00016",
309=>x"00016",
310=>x"00016",
311=>x"00016",
312=>x"00016",
313=>x"00016",
314=>x"00016",
315=>x"00016",
316=>x"00016",
317=>x"00016",
318=>x"00016",
319=>x"00016",
320=>x"00016",
321=>x"00016",
322=>x"00017",
323=>x"00017",
324=>x"00017",
325=>x"00017",
326=>x"00017",
327=>x"00017",
328=>x"00017",
329=>x"00017",
330=>x"00017",
331=>x"00017",
332=>x"00017",
333=>x"00017",
334=>x"00017",
335=>x"00017",
336=>x"00018",
337=>x"00018",
338=>x"00018",
339=>x"00018",
340=>x"00018",
341=>x"00018",
342=>x"00018",
343=>x"00018",
344=>x"00018",
345=>x"00018",
346=>x"00018",
347=>x"00018",
348=>x"00018",
349=>x"00018",
350=>x"00019",
351=>x"00019",
352=>x"00019",
353=>x"00019",
354=>x"00019",
355=>x"00019",
356=>x"00019",
357=>x"00019",
358=>x"00019",
359=>x"00019",
360=>x"00019",
361=>x"00019",
362=>x"00019",
363=>x"00019",
364=>x"0001a",
365=>x"0001a",
366=>x"0001a",
367=>x"0001a",
368=>x"0001a",
369=>x"0001a",
370=>x"0001a",
371=>x"0001a",
372=>x"0001a",
373=>x"0001a",
374=>x"0001a",
375=>x"0001a",
376=>x"0001a",
377=>x"0001a",
378=>x"0001b",
379=>x"0001b",
380=>x"0001b",
381=>x"0001b",
382=>x"0001b",
383=>x"0001b",
384=>x"0001b",
385=>x"0001b",
386=>x"0001b",
387=>x"0001b",
388=>x"0001b",
389=>x"0001b",
390=>x"0001b",
391=>x"0001b",
392=>x"0001c",
393=>x"0001c",
394=>x"0001c",
395=>x"0001c",
396=>x"0001c",
397=>x"0001c",
398=>x"0001c",
399=>x"0001c",
400=>x"0001c",
401=>x"0001c",
402=>x"0001c",
403=>x"0001c",
404=>x"0001c",
405=>x"0001c",
406=>x"0001d",
407=>x"0001d",
408=>x"0001d",
409=>x"0001d",
410=>x"0001d",
411=>x"0001d",
412=>x"0001d",
413=>x"0001d",
414=>x"0001d",
415=>x"0001d",
416=>x"0001d",
417=>x"0001d",
418=>x"0001d",
419=>x"0001d",
420=>x"0001e",
421=>x"0001e",
422=>x"0001e",
423=>x"0001e",
424=>x"0001e",
425=>x"0001e",
426=>x"0001e",
427=>x"0001e",
428=>x"0001e",
429=>x"0001e",
430=>x"0001e",
431=>x"0001e",
432=>x"0001e",
433=>x"0001e",
434=>x"0001f",
435=>x"0001f",
436=>x"0001f",
437=>x"0001f",
438=>x"0001f",
439=>x"0001f",
440=>x"0001f",
441=>x"0001f",
442=>x"0001f",
443=>x"0001f",
444=>x"0001f",
445=>x"0001f",
446=>x"0001f",
447=>x"0001f",
448=>x"00020",
449=>x"00020",
450=>x"00020",
451=>x"00020",
452=>x"00020",
453=>x"00020",
454=>x"00020",
455=>x"00020",
456=>x"00020",
457=>x"00020",
458=>x"00020",
459=>x"00020",
460=>x"00020",
461=>x"00020",
462=>x"00021",
463=>x"00021",
464=>x"00021",
465=>x"00021",
466=>x"00021",
467=>x"00021",
468=>x"00021",
469=>x"00021",
470=>x"00021",
471=>x"00021",
472=>x"00021",
473=>x"00021",
474=>x"00021",
475=>x"00021",
476=>x"00022",
477=>x"00022",
478=>x"00022",
479=>x"00022",
480=>x"00022",
481=>x"00022",
482=>x"00022",
483=>x"00022",
484=>x"00022",
485=>x"00022",
486=>x"00022",
487=>x"00022",
488=>x"00022",
489=>x"00022",
490=>x"00023",
491=>x"00023",
492=>x"00023",
493=>x"00023",
494=>x"00023",
495=>x"00023",
496=>x"00023",
497=>x"00023",
498=>x"00023",
499=>x"00023",
500=>x"00023",
501=>x"00023",
502=>x"00023",
503=>x"00023",
504=>x"00024",
505=>x"00024",
506=>x"00024",
507=>x"00024",
508=>x"00024",
509=>x"00024",
510=>x"00024",
511=>x"00024",
512=>x"00024",
513=>x"00024",
514=>x"00024",
515=>x"00024",
516=>x"00024",
517=>x"00024",
518=>x"00025",
519=>x"00025",
520=>x"00025",
521=>x"00025",
522=>x"00025",
523=>x"00025",
524=>x"00025",
525=>x"00025",
526=>x"00025",
527=>x"00025",
528=>x"00025",
529=>x"00025",
530=>x"00025",
531=>x"00025",
532=>x"00026",
533=>x"00026",
534=>x"00026",
535=>x"00026",
536=>x"00026",
537=>x"00026",
538=>x"00026",
539=>x"00026",
540=>x"00026",
541=>x"00026",
542=>x"00026",
543=>x"00026",
544=>x"00026",
545=>x"00026",
546=>x"00027",
547=>x"00027",
548=>x"00027",
549=>x"00027",
550=>x"00027",
551=>x"00027",
552=>x"00027",
553=>x"00027",
554=>x"00027",
555=>x"00027",
556=>x"00027",
557=>x"00027",
558=>x"00027",
559=>x"00027",
560=>x"00028",
561=>x"00028",
562=>x"00028",
563=>x"00028",
564=>x"00028",
565=>x"00028",
566=>x"00028",
567=>x"00028",
568=>x"00028",
569=>x"00028",
570=>x"00028",
571=>x"00028",
572=>x"00028",
573=>x"00028",
574=>x"00029",
575=>x"00029",
576=>x"00029",
577=>x"00029",
578=>x"00029",
579=>x"00029",
580=>x"00029",
581=>x"00029",
582=>x"00029",
583=>x"00029",
584=>x"00029",
585=>x"00029",
586=>x"00029",
587=>x"00029",
588=>x"0002a",
589=>x"0002a",
590=>x"0002a",
591=>x"0002a",
592=>x"0002a",
593=>x"0002a",
594=>x"0002a",
595=>x"0002a",
596=>x"0002a",
597=>x"0002a",
598=>x"0002a",
599=>x"0002a",
600=>x"0002a",
601=>x"0002a",
602=>x"0002b",
603=>x"0002b",
604=>x"0002b",
605=>x"0002b",
606=>x"0002b",
607=>x"0002b",
608=>x"0002b",
609=>x"0002b",
610=>x"0002b",
611=>x"0002b",
612=>x"0002b",
613=>x"0002b",
614=>x"0002b",
615=>x"0002b",
616=>x"0002c",
617=>x"0002c",
618=>x"0002c",
619=>x"0002c",
620=>x"0002c",
621=>x"0002c",
622=>x"0002c",
623=>x"0002c",
624=>x"0002c",
625=>x"0002c",
626=>x"0002c",
627=>x"0002c",
628=>x"0002c",
629=>x"0002c",
630=>x"0002d",
631=>x"0002d",
632=>x"0002d",
633=>x"0002d",
634=>x"0002d",
635=>x"0002d",
636=>x"0002d",
637=>x"0002d",
638=>x"0002d",
639=>x"0002d",
640=>x"0002d",
641=>x"0002d",
642=>x"0002d",
643=>x"0002d",
644=>x"0002e",
645=>x"0002e",
646=>x"0002e",
647=>x"0002e",
648=>x"0002e",
649=>x"0002e",
650=>x"0002e",
651=>x"0002e",
652=>x"0002e",
653=>x"0002e",
654=>x"0002e",
655=>x"0002e",
656=>x"0002e",
657=>x"0002e",
658=>x"0002f",
659=>x"0002f",
660=>x"0002f",
661=>x"0002f",
662=>x"0002f",
663=>x"0002f",
664=>x"0002f",
665=>x"0002f",
666=>x"0002f",
667=>x"0002f",
668=>x"0002f",
669=>x"0002f",
670=>x"0002f",
671=>x"0002f",
672=>x"00030",
673=>x"00030",
674=>x"00030",
675=>x"00030",
676=>x"00030",
677=>x"00030",
678=>x"00030",
679=>x"00030",
680=>x"00030",
681=>x"00030",
682=>x"00030",
683=>x"00030",
684=>x"00030",
685=>x"00030",
686=>x"00031",
687=>x"00031",
688=>x"00031",
689=>x"00031",
690=>x"00031",
691=>x"00031",
692=>x"00031",
693=>x"00031",
694=>x"00031",
695=>x"00031",
696=>x"00031",
697=>x"00031",
698=>x"00031",
699=>x"00031",
700=>x"00032",
701=>x"00032",
702=>x"00032",
703=>x"00032",
704=>x"00032",
705=>x"00032",
706=>x"00032",
707=>x"00032",
708=>x"00032",
709=>x"00032",
710=>x"00032",
711=>x"00032",
712=>x"00032",
713=>x"00032",
714=>x"00033",
715=>x"00033",
716=>x"00033",
717=>x"00033",
718=>x"00033",
719=>x"00033",
720=>x"00033",
721=>x"00033",
722=>x"00033",
723=>x"00033",
724=>x"00033",
725=>x"00033",
726=>x"00033",
727=>x"00033",
728=>x"00034",
729=>x"00034",
730=>x"00034",
731=>x"00034",
732=>x"00034",
733=>x"00034",
734=>x"00034",
735=>x"00034",
736=>x"00034",
737=>x"00034",
738=>x"00034",
739=>x"00034",
740=>x"00034",
741=>x"00034",
742=>x"00035",
743=>x"00035",
744=>x"00035",
745=>x"00035",
746=>x"00035",
747=>x"00035",
748=>x"00035",
749=>x"00035",
750=>x"00035",
751=>x"00035",
752=>x"00035",
753=>x"00035",
754=>x"00035",
755=>x"00035",
756=>x"00036",
757=>x"00036",
758=>x"00036",
759=>x"00036",
760=>x"00036",
761=>x"00036",
762=>x"00036",
763=>x"00036",
764=>x"00036",
765=>x"00036",
766=>x"00036",
767=>x"00036",
768=>x"00036",
769=>x"00036",
770=>x"00037",
771=>x"00037",
772=>x"00037",
773=>x"00037",
774=>x"00037",
775=>x"00037",
776=>x"00037",
777=>x"00037",
778=>x"00037",
779=>x"00037",
780=>x"00037",
781=>x"00037",
782=>x"00037",
783=>x"00037",
784=>x"00038",
785=>x"00038",
786=>x"00038",
787=>x"00038",
788=>x"00038",
789=>x"00038",
790=>x"00038",
791=>x"00038",
792=>x"00038",
793=>x"00038",
794=>x"00038",
795=>x"00038",
796=>x"00038",
797=>x"00038",
798=>x"00039",
799=>x"00039",
800=>x"00039",
801=>x"00039",
802=>x"00039",
803=>x"00039",
804=>x"00039",
805=>x"00039",
806=>x"00039",
807=>x"00039",
808=>x"00039",
809=>x"00039",
810=>x"00039",
811=>x"00039",
812=>x"0003a",
813=>x"0003a",
814=>x"0003a",
815=>x"0003a",
816=>x"0003a",
817=>x"0003a",
818=>x"0003a",
819=>x"0003a",
820=>x"0003a",
821=>x"0003a",
822=>x"0003a",
823=>x"0003a",
824=>x"0003a",
825=>x"0003a",
826=>x"0003b",
827=>x"0003b",
828=>x"0003b",
829=>x"0003b",
830=>x"0003b",
831=>x"0003b",
832=>x"0003b",
833=>x"0003b",
834=>x"0003b",
835=>x"0003b",
836=>x"0003b",
837=>x"0003b",
838=>x"0003b",
839=>x"0003b",
840=>x"0003c",
841=>x"0003c",
842=>x"0003c",
843=>x"0003c",
844=>x"0003c",
845=>x"0003c",
846=>x"0003c",
847=>x"0003c",
848=>x"0003c",
849=>x"0003c",
850=>x"0003c",
851=>x"0003c",
852=>x"0003c",
853=>x"0003c",
854=>x"0003d",
855=>x"0003d",
856=>x"0003d",
857=>x"0003d",
858=>x"0003d",
859=>x"0003d",
860=>x"0003d",
861=>x"0003d",
862=>x"0003d",
863=>x"0003d",
864=>x"0003d",
865=>x"0003d",
866=>x"0003d",
867=>x"0003d",
868=>x"0003e",
869=>x"0003e",
870=>x"0003e",
871=>x"0003e",
872=>x"0003e",
873=>x"0003e",
874=>x"0003e",
875=>x"0003e",
876=>x"0003e",
877=>x"0003e",
878=>x"0003e",
879=>x"0003e",
880=>x"0003e",
881=>x"0003e",
882=>x"0003f",
883=>x"0003f",
884=>x"0003f",
885=>x"0003f",
886=>x"0003f",
887=>x"0003f",
888=>x"0003f",
889=>x"0003f",
890=>x"0003f",
891=>x"0003f",
892=>x"0003f",
893=>x"0003f",
894=>x"0003f",
895=>x"0003f",
896=>x"00040",
897=>x"00040",
898=>x"00040",
899=>x"00040",
900=>x"00040",
901=>x"00040",
902=>x"00040",
903=>x"00040",
904=>x"00040",
905=>x"00040",
906=>x"00040",
907=>x"00040",
908=>x"00040",
909=>x"00040",
910=>x"00041",
911=>x"00041",
912=>x"00041",
913=>x"00041",
914=>x"00041",
915=>x"00041",
916=>x"00041",
917=>x"00041",
918=>x"00041",
919=>x"00041",
920=>x"00041",
921=>x"00041",
922=>x"00041",
923=>x"00041",
924=>x"00042",
925=>x"00042",
926=>x"00042",
927=>x"00042",
928=>x"00042",
929=>x"00042",
930=>x"00042",
931=>x"00042",
932=>x"00042",
933=>x"00042",
934=>x"00042",
935=>x"00042",
936=>x"00042",
937=>x"00042",
938=>x"00043",
939=>x"00043",
940=>x"00043",
941=>x"00043",
942=>x"00043",
943=>x"00043",
944=>x"00043",
945=>x"00043",
946=>x"00043",
947=>x"00043",
948=>x"00043",
949=>x"00043",
950=>x"00043",
951=>x"00043",
952=>x"00044",
953=>x"00044",
954=>x"00044",
955=>x"00044",
956=>x"00044",
957=>x"00044",
958=>x"00044",
959=>x"00044",
960=>x"00044",
961=>x"00044",
962=>x"00044",
963=>x"00044",
964=>x"00044",
965=>x"00044",
966=>x"00045",
967=>x"00045",
968=>x"00045",
969=>x"00045",
970=>x"00045",
971=>x"00045",
972=>x"00045",
973=>x"00045",
974=>x"00045",
975=>x"00045",
976=>x"00045",
977=>x"00045",
978=>x"00045",
979=>x"00045",
980=>x"00046",
981=>x"00046",
982=>x"00046",
983=>x"00046",
984=>x"00046",
985=>x"00046",
986=>x"00046",
987=>x"00046",
988=>x"00046",
989=>x"00046",
990=>x"00046",
991=>x"00046",
992=>x"00046",
993=>x"00046",
994=>x"00047",
995=>x"00047",
996=>x"00047",
997=>x"00047",
998=>x"00047",
999=>x"00047",
1000=>x"00047",
1001=>x"00047",
1002=>x"00047",
1003=>x"00047",
1004=>x"00047",
1005=>x"00047",
1006=>x"00047",
1007=>x"00047",
1008=>x"00048",
1009=>x"00048",
1010=>x"00048",
1011=>x"00048",
1012=>x"00048",
1013=>x"00048",
1014=>x"00048",
1015=>x"00048",
1016=>x"00048",
1017=>x"00048",
1018=>x"00048",
1019=>x"00048",
1020=>x"00048",
1021=>x"00048",
1022=>x"00049",
1023=>x"00049",
1024=>x"00049",
1025=>x"00049",
1026=>x"00049",
1027=>x"00049",
1028=>x"00049",
1029=>x"00049",
1030=>x"00049",
1031=>x"00049",
1032=>x"00049",
1033=>x"00049",
1034=>x"00049",
1035=>x"00049",
1036=>x"0004a",
1037=>x"0004a",
1038=>x"0004a",
1039=>x"0004a",
1040=>x"0004a",
1041=>x"0004a",
1042=>x"0004a",
1043=>x"0004a",
1044=>x"0004a",
1045=>x"0004a",
1046=>x"0004a",
1047=>x"0004a",
1048=>x"0004a",
1049=>x"0004a",
1050=>x"0004b",
1051=>x"0004b",
1052=>x"0004b",
1053=>x"0004b",
1054=>x"0004b",
1055=>x"0004b",
1056=>x"0004b",
1057=>x"0004b",
1058=>x"0004b",
1059=>x"0004b",
1060=>x"0004b",
1061=>x"0004b",
1062=>x"0004b",
1063=>x"0004b",
1064=>x"0004c",
1065=>x"0004c",
1066=>x"0004c",
1067=>x"0004c",
1068=>x"0004c",
1069=>x"0004c",
1070=>x"0004c",
1071=>x"0004c",
1072=>x"0004c",
1073=>x"0004c",
1074=>x"0004c",
1075=>x"0004c",
1076=>x"0004c",
1077=>x"0004c",
1078=>x"0004d",
1079=>x"0004d",
1080=>x"0004d",
1081=>x"0004d",
1082=>x"0004d",
1083=>x"0004d",
1084=>x"0004d",
1085=>x"0004d",
1086=>x"0004d",
1087=>x"0004d",
1088=>x"0004d",
1089=>x"0004d",
1090=>x"0004d",
1091=>x"0004d",
1092=>x"0004e",
1093=>x"0004e",
1094=>x"0004e",
1095=>x"0004e",
1096=>x"0004e",
1097=>x"0004e",
1098=>x"0004e",
1099=>x"0004e",
1100=>x"0004e",
1101=>x"0004e",
1102=>x"0004e",
1103=>x"0004e",
1104=>x"0004e",
1105=>x"0004e",
1106=>x"0004f",
1107=>x"0004f",
1108=>x"0004f",
1109=>x"0004f",
1110=>x"0004f",
1111=>x"0004f",
1112=>x"0004f",
1113=>x"0004f",
1114=>x"0004f",
1115=>x"0004f",
1116=>x"0004f",
1117=>x"0004f",
1118=>x"0004f",
1119=>x"0004f",
1120=>x"00050",
1121=>x"00050",
1122=>x"00050",
1123=>x"00050",
1124=>x"00050",
1125=>x"00050",
1126=>x"00050",
1127=>x"00050",
1128=>x"00050",
1129=>x"00050",
1130=>x"00050",
1131=>x"00050",
1132=>x"00050",
1133=>x"00050",
1134=>x"00051",
1135=>x"00051",
1136=>x"00051",
1137=>x"00051",
1138=>x"00051",
1139=>x"00051",
1140=>x"00051",
1141=>x"00051",
1142=>x"00051",
1143=>x"00051",
1144=>x"00051",
1145=>x"00051",
1146=>x"00051",
1147=>x"00051",
1148=>x"00052",
1149=>x"00052",
1150=>x"00052",
1151=>x"00052",
1152=>x"00052",
1153=>x"00052",
1154=>x"00052",
1155=>x"00052",
1156=>x"00052",
1157=>x"00052",
1158=>x"00052",
1159=>x"00052",
1160=>x"00052",
1161=>x"00052",
1162=>x"00053",
1163=>x"00053",
1164=>x"00053",
1165=>x"00053",
1166=>x"00053",
1167=>x"00053",
1168=>x"00053",
1169=>x"00053",
1170=>x"00053",
1171=>x"00053",
1172=>x"00053",
1173=>x"00053",
1174=>x"00053",
1175=>x"00053",
1176=>x"00054",
1177=>x"00054",
1178=>x"00054",
1179=>x"00054",
1180=>x"00054",
1181=>x"00054",
1182=>x"00054",
1183=>x"00054",
1184=>x"00054",
1185=>x"00054",
1186=>x"00054",
1187=>x"00054",
1188=>x"00054",
1189=>x"00054",
1190=>x"00055",
1191=>x"00055",
1192=>x"00055",
1193=>x"00055",
1194=>x"00055",
1195=>x"00055",
1196=>x"00055",
1197=>x"00055",
1198=>x"00055",
1199=>x"00055",
1200=>x"00055",
1201=>x"00055",
1202=>x"00055",
1203=>x"00055",
1204=>x"00056",
1205=>x"00056",
1206=>x"00056",
1207=>x"00056",
1208=>x"00056",
1209=>x"00056",
1210=>x"00056",
1211=>x"00056",
1212=>x"00056",
1213=>x"00056",
1214=>x"00056",
1215=>x"00056",
1216=>x"00056",
1217=>x"00056",
1218=>x"00057",
1219=>x"00057",
1220=>x"00057",
1221=>x"00057",
1222=>x"00057",
1223=>x"00057",
1224=>x"00057",
1225=>x"00057",
1226=>x"00057",
1227=>x"00057",
1228=>x"00057",
1229=>x"00057",
1230=>x"00057",
1231=>x"00057",
1232=>x"00058",
1233=>x"00058",
1234=>x"00058",
1235=>x"00058",
1236=>x"00058",
1237=>x"00058",
1238=>x"00058",
1239=>x"00058",
1240=>x"00058",
1241=>x"00058",
1242=>x"00058",
1243=>x"00058",
1244=>x"00058",
1245=>x"00058",
1246=>x"00059",
1247=>x"00059",
1248=>x"00059",
1249=>x"00059",
1250=>x"00059",
1251=>x"00059",
1252=>x"00059",
1253=>x"00059",
1254=>x"00059",
1255=>x"00059",
1256=>x"00059",
1257=>x"00059",
1258=>x"00059",
1259=>x"00059",
1260=>x"0005a",
1261=>x"0005a",
1262=>x"0005a",
1263=>x"0005a",
1264=>x"0005a",
1265=>x"0005a",
1266=>x"0005a",
1267=>x"0005a",
1268=>x"0005a",
1269=>x"0005a",
1270=>x"0005a",
1271=>x"0005a",
1272=>x"0005a",
1273=>x"0005a",
1274=>x"0005b",
1275=>x"0005b",
1276=>x"0005b",
1277=>x"0005b",
1278=>x"0005b",
1279=>x"0005b",
1280=>x"0005b",
1281=>x"0005b",
1282=>x"0005b",
1283=>x"0005b",
1284=>x"0005b",
1285=>x"0005b",
1286=>x"0005b",
1287=>x"0005b",
1288=>x"0005c",
1289=>x"0005c",
1290=>x"0005c",
1291=>x"0005c",
1292=>x"0005c",
1293=>x"0005c",
1294=>x"0005c",
1295=>x"0005c",
1296=>x"0005c",
1297=>x"0005c",
1298=>x"0005c",
1299=>x"0005c",
1300=>x"0005c",
1301=>x"0005c",
1302=>x"0005d",
1303=>x"0005d",
1304=>x"0005d",
1305=>x"0005d",
1306=>x"0005d",
1307=>x"0005d",
1308=>x"0005d",
1309=>x"0005d",
1310=>x"0005d",
1311=>x"0005d",
1312=>x"0005d",
1313=>x"0005d",
1314=>x"0005d",
1315=>x"0005d",
1316=>x"0005e",
1317=>x"0005e",
1318=>x"0005e",
1319=>x"0005e",
1320=>x"0005e",
1321=>x"0005e",
1322=>x"0005e",
1323=>x"0005e",
1324=>x"0005e",
1325=>x"0005e",
1326=>x"0005e",
1327=>x"0005e",
1328=>x"0005e",
1329=>x"0005e",
1330=>x"0005f",
1331=>x"0005f",
1332=>x"0005f",
1333=>x"0005f",
1334=>x"0005f",
1335=>x"0005f",
1336=>x"0005f",
1337=>x"0005f",
1338=>x"0005f",
1339=>x"0005f",
1340=>x"0005f",
1341=>x"0005f",
1342=>x"0005f",
1343=>x"0005f",
1344=>x"00060",
1345=>x"00060",
1346=>x"00060",
1347=>x"00060",
1348=>x"00060",
1349=>x"00060",
1350=>x"00060",
1351=>x"00060",
1352=>x"00060",
1353=>x"00060",
1354=>x"00060",
1355=>x"00060",
1356=>x"00060",
1357=>x"00060",
1358=>x"00061",
1359=>x"00061",
1360=>x"00061",
1361=>x"00061",
1362=>x"00061",
1363=>x"00061",
1364=>x"00061",
1365=>x"00061",
1366=>x"00061",
1367=>x"00061",
1368=>x"00061",
1369=>x"00061",
1370=>x"00061",
1371=>x"00061",
1372=>x"00062",
1373=>x"00062",
1374=>x"00062",
1375=>x"00062",
1376=>x"00062",
1377=>x"00062",
1378=>x"00062",
1379=>x"00062",
1380=>x"00062",
1381=>x"00062",
1382=>x"00062",
1383=>x"00062",
1384=>x"00062",
1385=>x"00062",
1386=>x"00063",
1387=>x"00063",
1388=>x"00063",
1389=>x"00063",
1390=>x"00063",
1391=>x"00063",
1392=>x"00063",
1393=>x"00063",
1394=>x"00063",
1395=>x"00063",
1396=>x"00063",
1397=>x"00063",
1398=>x"00063",
1399=>x"00063",
1400=>x"00064"
);
begin
Cout<=memory(to_integer(unsigned(addr)));

end Behavioral;
